LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE ALUPaket IS

COMPONENT arit_jedinica IS
	PORT (Ulaz1, Ulaz2:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
			Izlaz			:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			Selekcija	:	IN  STD_LOGIC_VECTOR(2 DOWNTO 0)
		);
END COMPONENT;

COMPONENT log_jedinica IS
	PORT( Ulaz1, Ulaz2	:	IN    STD_LOGIC_VECTOR(7 DOWNTO 0);
			Izlaz				: 	OUT	STD_LOGIC_VECTOR(7 DOWNTO 0);
			Selekcija		:	IN		STD_LOGIC_VECTOR(2 DOWNTO 0)
			);
END COMPONENT;

COMPONENT multipleksor IS

			PORT(
			Ulaz1, Ulaz2:	IN	 STD_LOGIC_VECTOR(7 DOWNTO 0);
			Izlaz			:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			Selekcija	:	IN	 STD_LOGIC
	);
	
END COMPONENT;

END PACKAGE ALUPaket;